`timescale 1ns / 1ps


module tb_mux_8to1(

    );
    
    reg a0, a1, a2, a3, a4, a5, a6, a7;
    reg s0, s1, s2;
    
    wire y;
    
    mux_8to1 uut(a0, a1, a2, a3, a4, a5, a6,a7, s0, s1, s2, y);
    
    initial begin
    
    s0 = 0; s1 = 0; s2 = 0; //000
    a0 = 1; a1 = 0; a2 = 0; a3 = 0; a4 = 0; a5 = 0; a6 = 0; a7 = 0;
    #10; // a0
    
    s0 = 0; s1 = 0; s2 = 1; // 001
    a0 = 0; a1 = 1; a2 = 0; a3 = 0; a4 = 0; a5 = 0; a6 = 0; a7 = 0;
    #10; //a
    
    s0 = 0; s1 = 1; s2 = 0; //010 
    a0 = 0; a1 = 0; a2 = 1; a3 = 0; a4 = 0; a5 = 0; a6 = 0; a7 = 0;
    #10; // a2
    
    s0 = 0; s1 = 1; s2 = 1;// 011
    a0 = 0; a1 = 0; a2 = 0; a3 = 1; a4 = 0; a5 = 0; a6 = 0; a7 = 0;
    #10; //a3
    
    s0 = 1; s1 = 0; s2 = 0; //100
    a0 = 0; a1 = 0; a2 = 0; a3 = 0; a4 = 1; a5 = 0; a6 = 0; a7 = 0;
    #10; //a4
    
    s0 = 1; s1 = 0; s2 = 1; //101
    a0 = 0; a1 = 0; a2 = 0; a3 = 0; a4 = 0; a5 = 1; a6 = 0; a7 = 0;
    #10; //a5
    
    s0 = 1; s1 = 1; s2 = 0; //110
    a0 = 0; a1 = 0; a2 = 0; a3 = 0; a4 = 0; a5 = 0; a6 = 1; a7 = 0;
    #10; //a6
    
    s0 = 1; s1 = 1; s2 = 1; //111
    a0 = 0; a1 = 0; a2 = 0; a3 = 0; a4 = 0; a5 = 0; a6 = 0; a7 = 1;
    //a7
    
    $finish;
    
    end
endmodule
