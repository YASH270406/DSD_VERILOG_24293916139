`timescale 1ns / 1ps

module tb_and_gate(

    );
    
reg a,b;
wire y;

and_gate uut(a, b, y);

initial begin

a = 0; b = 0;
#10;

a = 0; b = 1;
#10;

a = 1; b = 0;
#10;

a = 1; b = 1;

$finish;

end
endmodule
