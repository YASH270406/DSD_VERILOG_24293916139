`timescale 1ns / 1ps

module mux_4to1(

    input a, b, c, d, s0, s1,
    
    output y

    );
    
    assign y = ((~s0)&(~s1)&a) | ((~s0)&(s1)&b) 
    |((s0)&(~s1)&c) | ((s0)&(s1)&d);
endmodule
